// my_sys.v

// Generated using ACDS version 23.3 104

`timescale 1 ps / 1 ps
module my_sys (
		input  wire  clk_clk,     //   clk.clk
		input  wire  reset_reset  // reset.reset
	);

	wire         clock_in_out_clk_clk;                                 // clock_in:out_clk -> [mgc_axi4_master_0:ACLK, mm_interconnect_0:clock_in_out_clk_clk, my_sys_onchip_memory:clk, reset_in:clk, rst_controller:clk, rst_controller_001:clk]
	wire   [7:0] mgc_axi4_master_0_altera_axi4_master_ruser;           // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_ruser -> mgc_axi4_master_0:RUSER
	wire   [7:0] mgc_axi4_master_0_altera_axi4_master_wuser;           // mgc_axi4_master_0:WUSER -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wuser
	wire   [1:0] mgc_axi4_master_0_altera_axi4_master_awburst;         // mgc_axi4_master_0:AWBURST -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awburst
	wire   [3:0] mgc_axi4_master_0_altera_axi4_master_arregion;        // mgc_axi4_master_0:ARREGION -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arregion
	wire   [7:0] mgc_axi4_master_0_altera_axi4_master_arlen;           // mgc_axi4_master_0:ARLEN -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arlen
	wire   [3:0] mgc_axi4_master_0_altera_axi4_master_arqos;           // mgc_axi4_master_0:ARQOS -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arqos
	wire   [7:0] mgc_axi4_master_0_altera_axi4_master_awuser;          // mgc_axi4_master_0:AWUSER -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awuser
	wire         mgc_axi4_master_0_altera_axi4_master_wready;          // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wready -> mgc_axi4_master_0:WREADY
	wire   [3:0] mgc_axi4_master_0_altera_axi4_master_wstrb;           // mgc_axi4_master_0:WSTRB -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wstrb
	wire  [17:0] mgc_axi4_master_0_altera_axi4_master_rid;             // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rid -> mgc_axi4_master_0:RID
	wire         mgc_axi4_master_0_altera_axi4_master_rready;          // mgc_axi4_master_0:RREADY -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rready
	wire   [7:0] mgc_axi4_master_0_altera_axi4_master_awlen;           // mgc_axi4_master_0:AWLEN -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awlen
	wire   [3:0] mgc_axi4_master_0_altera_axi4_master_awqos;           // mgc_axi4_master_0:AWQOS -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awqos
	wire   [3:0] mgc_axi4_master_0_altera_axi4_master_arcache;         // mgc_axi4_master_0:ARCACHE -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arcache
	wire         mgc_axi4_master_0_altera_axi4_master_wvalid;          // mgc_axi4_master_0:WVALID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wvalid
	wire  [15:0] mgc_axi4_master_0_altera_axi4_master_araddr;          // mgc_axi4_master_0:ARADDR -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_araddr
	wire   [2:0] mgc_axi4_master_0_altera_axi4_master_arprot;          // mgc_axi4_master_0:ARPROT -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arprot
	wire   [2:0] mgc_axi4_master_0_altera_axi4_master_awprot;          // mgc_axi4_master_0:AWPROT -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awprot
	wire         mgc_axi4_master_0_altera_axi4_master_arvalid;         // mgc_axi4_master_0:ARVALID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arvalid
	wire  [31:0] mgc_axi4_master_0_altera_axi4_master_wdata;           // mgc_axi4_master_0:WDATA -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wdata
	wire   [3:0] mgc_axi4_master_0_altera_axi4_master_awcache;         // mgc_axi4_master_0:AWCACHE -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awcache
	wire  [17:0] mgc_axi4_master_0_altera_axi4_master_arid;            // mgc_axi4_master_0:ARID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arid
	wire         mgc_axi4_master_0_altera_axi4_master_arlock;          // mgc_axi4_master_0:ARLOCK -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arlock
	wire         mgc_axi4_master_0_altera_axi4_master_awlock;          // mgc_axi4_master_0:AWLOCK -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awlock
	wire  [15:0] mgc_axi4_master_0_altera_axi4_master_awaddr;          // mgc_axi4_master_0:AWADDR -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awaddr
	wire         mgc_axi4_master_0_altera_axi4_master_arready;         // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arready -> mgc_axi4_master_0:ARREADY
	wire   [1:0] mgc_axi4_master_0_altera_axi4_master_bresp;           // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_bresp -> mgc_axi4_master_0:BRESP
	wire  [31:0] mgc_axi4_master_0_altera_axi4_master_rdata;           // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rdata -> mgc_axi4_master_0:RDATA
	wire         mgc_axi4_master_0_altera_axi4_master_awready;         // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awready -> mgc_axi4_master_0:AWREADY
	wire   [1:0] mgc_axi4_master_0_altera_axi4_master_arburst;         // mgc_axi4_master_0:ARBURST -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arburst
	wire   [2:0] mgc_axi4_master_0_altera_axi4_master_arsize;          // mgc_axi4_master_0:ARSIZE -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arsize
	wire         mgc_axi4_master_0_altera_axi4_master_rlast;           // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rlast -> mgc_axi4_master_0:RLAST
	wire         mgc_axi4_master_0_altera_axi4_master_bready;          // mgc_axi4_master_0:BREADY -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_bready
	wire         mgc_axi4_master_0_altera_axi4_master_wlast;           // mgc_axi4_master_0:WLAST -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wlast
	wire   [3:0] mgc_axi4_master_0_altera_axi4_master_awregion;        // mgc_axi4_master_0:AWREGION -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awregion
	wire   [7:0] mgc_axi4_master_0_altera_axi4_master_buser;           // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_buser -> mgc_axi4_master_0:BUSER
	wire   [1:0] mgc_axi4_master_0_altera_axi4_master_rresp;           // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rresp -> mgc_axi4_master_0:RRESP
	wire  [17:0] mgc_axi4_master_0_altera_axi4_master_awid;            // mgc_axi4_master_0:AWID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awid
	wire  [17:0] mgc_axi4_master_0_altera_axi4_master_bid;             // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_bid -> mgc_axi4_master_0:BID
	wire         mgc_axi4_master_0_altera_axi4_master_bvalid;          // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_bvalid -> mgc_axi4_master_0:BVALID
	wire         mgc_axi4_master_0_altera_axi4_master_awvalid;         // mgc_axi4_master_0:AWVALID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awvalid
	wire   [2:0] mgc_axi4_master_0_altera_axi4_master_awsize;          // mgc_axi4_master_0:AWSIZE -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awsize
	wire         mgc_axi4_master_0_altera_axi4_master_rvalid;          // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rvalid -> mgc_axi4_master_0:RVALID
	wire   [7:0] mgc_axi4_master_0_altera_axi4_master_aruser;          // mgc_axi4_master_0:ARUSER -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_aruser
	wire         mm_interconnect_0_my_sys_onchip_memory_s1_chipselect; // mm_interconnect_0:my_sys_onchip_memory_s1_chipselect -> my_sys_onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_my_sys_onchip_memory_s1_readdata;   // my_sys_onchip_memory:readdata -> mm_interconnect_0:my_sys_onchip_memory_s1_readdata
	wire   [6:0] mm_interconnect_0_my_sys_onchip_memory_s1_address;    // mm_interconnect_0:my_sys_onchip_memory_s1_address -> my_sys_onchip_memory:address
	wire   [3:0] mm_interconnect_0_my_sys_onchip_memory_s1_byteenable; // mm_interconnect_0:my_sys_onchip_memory_s1_byteenable -> my_sys_onchip_memory:byteenable
	wire         mm_interconnect_0_my_sys_onchip_memory_s1_write;      // mm_interconnect_0:my_sys_onchip_memory_s1_write -> my_sys_onchip_memory:write
	wire  [31:0] mm_interconnect_0_my_sys_onchip_memory_s1_writedata;  // mm_interconnect_0:my_sys_onchip_memory_s1_writedata -> my_sys_onchip_memory:writedata
	wire         mm_interconnect_0_my_sys_onchip_memory_s1_clken;      // mm_interconnect_0:my_sys_onchip_memory_s1_clken -> my_sys_onchip_memory:clken
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [mgc_axi4_master_0:ARESETn, my_sys_onchip_memory:reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> my_sys_onchip_memory:reset_req
	wire         reset_in_out_reset_reset;                             // reset_in:out_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                   // rst_controller_001:reset_out -> [mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mgc_axi4_master_0_reset_sink_reset_bridge_in_reset_reset]

	my_sys_clock_in clock_in (
		.in_clk  (clk_clk),              //   input,  width = 1,  in_clk.clk
		.out_clk (clock_in_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	my_sys_mgc_axi4_master_0 mgc_axi4_master_0 (
		.AWVALID  (mgc_axi4_master_0_altera_axi4_master_awvalid),  //  output,   width = 1, altera_axi4_master.awvalid
		.AWPROT   (mgc_axi4_master_0_altera_axi4_master_awprot),   //  output,   width = 3,                   .awprot
		.AWREGION (mgc_axi4_master_0_altera_axi4_master_awregion), //  output,   width = 4,                   .awregion
		.AWLEN    (mgc_axi4_master_0_altera_axi4_master_awlen),    //  output,   width = 8,                   .awlen
		.AWSIZE   (mgc_axi4_master_0_altera_axi4_master_awsize),   //  output,   width = 3,                   .awsize
		.AWBURST  (mgc_axi4_master_0_altera_axi4_master_awburst),  //  output,   width = 2,                   .awburst
		.AWLOCK   (mgc_axi4_master_0_altera_axi4_master_awlock),   //  output,   width = 1,                   .awlock
		.AWCACHE  (mgc_axi4_master_0_altera_axi4_master_awcache),  //  output,   width = 4,                   .awcache
		.AWQOS    (mgc_axi4_master_0_altera_axi4_master_awqos),    //  output,   width = 4,                   .awqos
		.AWREADY  (mgc_axi4_master_0_altera_axi4_master_awready),  //   input,   width = 1,                   .awready
		.ARVALID  (mgc_axi4_master_0_altera_axi4_master_arvalid),  //  output,   width = 1,                   .arvalid
		.ARPROT   (mgc_axi4_master_0_altera_axi4_master_arprot),   //  output,   width = 3,                   .arprot
		.ARREGION (mgc_axi4_master_0_altera_axi4_master_arregion), //  output,   width = 4,                   .arregion
		.ARLEN    (mgc_axi4_master_0_altera_axi4_master_arlen),    //  output,   width = 8,                   .arlen
		.ARSIZE   (mgc_axi4_master_0_altera_axi4_master_arsize),   //  output,   width = 3,                   .arsize
		.ARBURST  (mgc_axi4_master_0_altera_axi4_master_arburst),  //  output,   width = 2,                   .arburst
		.ARLOCK   (mgc_axi4_master_0_altera_axi4_master_arlock),   //  output,   width = 1,                   .arlock
		.ARCACHE  (mgc_axi4_master_0_altera_axi4_master_arcache),  //  output,   width = 4,                   .arcache
		.ARQOS    (mgc_axi4_master_0_altera_axi4_master_arqos),    //  output,   width = 4,                   .arqos
		.ARREADY  (mgc_axi4_master_0_altera_axi4_master_arready),  //   input,   width = 1,                   .arready
		.RVALID   (mgc_axi4_master_0_altera_axi4_master_rvalid),   //   input,   width = 1,                   .rvalid
		.RRESP    (mgc_axi4_master_0_altera_axi4_master_rresp),    //   input,   width = 2,                   .rresp
		.RLAST    (mgc_axi4_master_0_altera_axi4_master_rlast),    //   input,   width = 1,                   .rlast
		.RREADY   (mgc_axi4_master_0_altera_axi4_master_rready),   //  output,   width = 1,                   .rready
		.WVALID   (mgc_axi4_master_0_altera_axi4_master_wvalid),   //  output,   width = 1,                   .wvalid
		.WLAST    (mgc_axi4_master_0_altera_axi4_master_wlast),    //  output,   width = 1,                   .wlast
		.WREADY   (mgc_axi4_master_0_altera_axi4_master_wready),   //   input,   width = 1,                   .wready
		.BVALID   (mgc_axi4_master_0_altera_axi4_master_bvalid),   //   input,   width = 1,                   .bvalid
		.BRESP    (mgc_axi4_master_0_altera_axi4_master_bresp),    //   input,   width = 2,                   .bresp
		.BREADY   (mgc_axi4_master_0_altera_axi4_master_bready),   //  output,   width = 1,                   .bready
		.AWADDR   (mgc_axi4_master_0_altera_axi4_master_awaddr),   //  output,  width = 16,                   .awaddr
		.AWID     (mgc_axi4_master_0_altera_axi4_master_awid),     //  output,  width = 18,                   .awid
		.AWUSER   (mgc_axi4_master_0_altera_axi4_master_awuser),   //  output,   width = 8,                   .awuser
		.ARADDR   (mgc_axi4_master_0_altera_axi4_master_araddr),   //  output,  width = 16,                   .araddr
		.ARID     (mgc_axi4_master_0_altera_axi4_master_arid),     //  output,  width = 18,                   .arid
		.ARUSER   (mgc_axi4_master_0_altera_axi4_master_aruser),   //  output,   width = 8,                   .aruser
		.RUSER    (mgc_axi4_master_0_altera_axi4_master_ruser),    //   input,   width = 8,                   .ruser
		.WUSER    (mgc_axi4_master_0_altera_axi4_master_wuser),    //  output,   width = 8,                   .wuser
		.BUSER    (mgc_axi4_master_0_altera_axi4_master_buser),    //   input,   width = 8,                   .buser
		.RDATA    (mgc_axi4_master_0_altera_axi4_master_rdata),    //   input,  width = 32,                   .rdata
		.RID      (mgc_axi4_master_0_altera_axi4_master_rid),      //   input,  width = 18,                   .rid
		.WDATA    (mgc_axi4_master_0_altera_axi4_master_wdata),    //  output,  width = 32,                   .wdata
		.WSTRB    (mgc_axi4_master_0_altera_axi4_master_wstrb),    //  output,   width = 4,                   .wstrb
		.BID      (mgc_axi4_master_0_altera_axi4_master_bid),      //   input,  width = 18,                   .bid
		.ACLK     (clock_in_out_clk_clk),                          //   input,   width = 1,         clock_sink.clk
		.ARESETn  (~rst_controller_reset_out_reset)                //   input,   width = 1,         reset_sink.reset_n
	);

	my_sys_onchip_memory my_sys_onchip_memory (
		.clk        (clock_in_out_clk_clk),                                 //   input,   width = 1,   clk1.clk
		.address    (mm_interconnect_0_my_sys_onchip_memory_s1_address),    //   input,   width = 7,     s1.address
		.clken      (mm_interconnect_0_my_sys_onchip_memory_s1_clken),      //   input,   width = 1,       .clken
		.chipselect (mm_interconnect_0_my_sys_onchip_memory_s1_chipselect), //   input,   width = 1,       .chipselect
		.write      (mm_interconnect_0_my_sys_onchip_memory_s1_write),      //   input,   width = 1,       .write
		.readdata   (mm_interconnect_0_my_sys_onchip_memory_s1_readdata),   //  output,  width = 32,       .readdata
		.writedata  (mm_interconnect_0_my_sys_onchip_memory_s1_writedata),  //   input,  width = 32,       .writedata
		.byteenable (mm_interconnect_0_my_sys_onchip_memory_s1_byteenable), //   input,   width = 4,       .byteenable
		.reset      (rst_controller_reset_out_reset),                       //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                    //   input,   width = 1,       .reset_req
	);

	my_sys_reset_in reset_in (
		.clk       (clock_in_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset  (reset_reset),              //   input,  width = 1,  in_reset.reset
		.out_reset (reset_in_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	my_sys_altera_mm_interconnect_1920_j74kjai mm_interconnect_0 (
		.mgc_axi4_master_0_altera_axi4_master_awid                                             (mgc_axi4_master_0_altera_axi4_master_awid),            //   input,  width = 18,                                            mgc_axi4_master_0_altera_axi4_master.awid
		.mgc_axi4_master_0_altera_axi4_master_awaddr                                           (mgc_axi4_master_0_altera_axi4_master_awaddr),          //   input,  width = 16,                                                                                .awaddr
		.mgc_axi4_master_0_altera_axi4_master_awlen                                            (mgc_axi4_master_0_altera_axi4_master_awlen),           //   input,   width = 8,                                                                                .awlen
		.mgc_axi4_master_0_altera_axi4_master_awsize                                           (mgc_axi4_master_0_altera_axi4_master_awsize),          //   input,   width = 3,                                                                                .awsize
		.mgc_axi4_master_0_altera_axi4_master_awburst                                          (mgc_axi4_master_0_altera_axi4_master_awburst),         //   input,   width = 2,                                                                                .awburst
		.mgc_axi4_master_0_altera_axi4_master_awlock                                           (mgc_axi4_master_0_altera_axi4_master_awlock),          //   input,   width = 1,                                                                                .awlock
		.mgc_axi4_master_0_altera_axi4_master_awcache                                          (mgc_axi4_master_0_altera_axi4_master_awcache),         //   input,   width = 4,                                                                                .awcache
		.mgc_axi4_master_0_altera_axi4_master_awprot                                           (mgc_axi4_master_0_altera_axi4_master_awprot),          //   input,   width = 3,                                                                                .awprot
		.mgc_axi4_master_0_altera_axi4_master_awuser                                           (mgc_axi4_master_0_altera_axi4_master_awuser),          //   input,   width = 8,                                                                                .awuser
		.mgc_axi4_master_0_altera_axi4_master_awqos                                            (mgc_axi4_master_0_altera_axi4_master_awqos),           //   input,   width = 4,                                                                                .awqos
		.mgc_axi4_master_0_altera_axi4_master_awregion                                         (mgc_axi4_master_0_altera_axi4_master_awregion),        //   input,   width = 4,                                                                                .awregion
		.mgc_axi4_master_0_altera_axi4_master_awvalid                                          (mgc_axi4_master_0_altera_axi4_master_awvalid),         //   input,   width = 1,                                                                                .awvalid
		.mgc_axi4_master_0_altera_axi4_master_awready                                          (mgc_axi4_master_0_altera_axi4_master_awready),         //  output,   width = 1,                                                                                .awready
		.mgc_axi4_master_0_altera_axi4_master_wdata                                            (mgc_axi4_master_0_altera_axi4_master_wdata),           //   input,  width = 32,                                                                                .wdata
		.mgc_axi4_master_0_altera_axi4_master_wstrb                                            (mgc_axi4_master_0_altera_axi4_master_wstrb),           //   input,   width = 4,                                                                                .wstrb
		.mgc_axi4_master_0_altera_axi4_master_wlast                                            (mgc_axi4_master_0_altera_axi4_master_wlast),           //   input,   width = 1,                                                                                .wlast
		.mgc_axi4_master_0_altera_axi4_master_wvalid                                           (mgc_axi4_master_0_altera_axi4_master_wvalid),          //   input,   width = 1,                                                                                .wvalid
		.mgc_axi4_master_0_altera_axi4_master_wuser                                            (mgc_axi4_master_0_altera_axi4_master_wuser),           //   input,   width = 8,                                                                                .wuser
		.mgc_axi4_master_0_altera_axi4_master_wready                                           (mgc_axi4_master_0_altera_axi4_master_wready),          //  output,   width = 1,                                                                                .wready
		.mgc_axi4_master_0_altera_axi4_master_bid                                              (mgc_axi4_master_0_altera_axi4_master_bid),             //  output,  width = 18,                                                                                .bid
		.mgc_axi4_master_0_altera_axi4_master_bresp                                            (mgc_axi4_master_0_altera_axi4_master_bresp),           //  output,   width = 2,                                                                                .bresp
		.mgc_axi4_master_0_altera_axi4_master_buser                                            (mgc_axi4_master_0_altera_axi4_master_buser),           //  output,   width = 8,                                                                                .buser
		.mgc_axi4_master_0_altera_axi4_master_bvalid                                           (mgc_axi4_master_0_altera_axi4_master_bvalid),          //  output,   width = 1,                                                                                .bvalid
		.mgc_axi4_master_0_altera_axi4_master_bready                                           (mgc_axi4_master_0_altera_axi4_master_bready),          //   input,   width = 1,                                                                                .bready
		.mgc_axi4_master_0_altera_axi4_master_arid                                             (mgc_axi4_master_0_altera_axi4_master_arid),            //   input,  width = 18,                                                                                .arid
		.mgc_axi4_master_0_altera_axi4_master_araddr                                           (mgc_axi4_master_0_altera_axi4_master_araddr),          //   input,  width = 16,                                                                                .araddr
		.mgc_axi4_master_0_altera_axi4_master_arlen                                            (mgc_axi4_master_0_altera_axi4_master_arlen),           //   input,   width = 8,                                                                                .arlen
		.mgc_axi4_master_0_altera_axi4_master_arsize                                           (mgc_axi4_master_0_altera_axi4_master_arsize),          //   input,   width = 3,                                                                                .arsize
		.mgc_axi4_master_0_altera_axi4_master_arburst                                          (mgc_axi4_master_0_altera_axi4_master_arburst),         //   input,   width = 2,                                                                                .arburst
		.mgc_axi4_master_0_altera_axi4_master_arlock                                           (mgc_axi4_master_0_altera_axi4_master_arlock),          //   input,   width = 1,                                                                                .arlock
		.mgc_axi4_master_0_altera_axi4_master_arcache                                          (mgc_axi4_master_0_altera_axi4_master_arcache),         //   input,   width = 4,                                                                                .arcache
		.mgc_axi4_master_0_altera_axi4_master_arprot                                           (mgc_axi4_master_0_altera_axi4_master_arprot),          //   input,   width = 3,                                                                                .arprot
		.mgc_axi4_master_0_altera_axi4_master_aruser                                           (mgc_axi4_master_0_altera_axi4_master_aruser),          //   input,   width = 8,                                                                                .aruser
		.mgc_axi4_master_0_altera_axi4_master_arqos                                            (mgc_axi4_master_0_altera_axi4_master_arqos),           //   input,   width = 4,                                                                                .arqos
		.mgc_axi4_master_0_altera_axi4_master_arregion                                         (mgc_axi4_master_0_altera_axi4_master_arregion),        //   input,   width = 4,                                                                                .arregion
		.mgc_axi4_master_0_altera_axi4_master_arvalid                                          (mgc_axi4_master_0_altera_axi4_master_arvalid),         //   input,   width = 1,                                                                                .arvalid
		.mgc_axi4_master_0_altera_axi4_master_arready                                          (mgc_axi4_master_0_altera_axi4_master_arready),         //  output,   width = 1,                                                                                .arready
		.mgc_axi4_master_0_altera_axi4_master_rid                                              (mgc_axi4_master_0_altera_axi4_master_rid),             //  output,  width = 18,                                                                                .rid
		.mgc_axi4_master_0_altera_axi4_master_rdata                                            (mgc_axi4_master_0_altera_axi4_master_rdata),           //  output,  width = 32,                                                                                .rdata
		.mgc_axi4_master_0_altera_axi4_master_rresp                                            (mgc_axi4_master_0_altera_axi4_master_rresp),           //  output,   width = 2,                                                                                .rresp
		.mgc_axi4_master_0_altera_axi4_master_rlast                                            (mgc_axi4_master_0_altera_axi4_master_rlast),           //  output,   width = 1,                                                                                .rlast
		.mgc_axi4_master_0_altera_axi4_master_rvalid                                           (mgc_axi4_master_0_altera_axi4_master_rvalid),          //  output,   width = 1,                                                                                .rvalid
		.mgc_axi4_master_0_altera_axi4_master_rready                                           (mgc_axi4_master_0_altera_axi4_master_rready),          //   input,   width = 1,                                                                                .rready
		.mgc_axi4_master_0_altera_axi4_master_ruser                                            (mgc_axi4_master_0_altera_axi4_master_ruser),           //  output,   width = 8,                                                                                .ruser
		.my_sys_onchip_memory_s1_address                                                       (mm_interconnect_0_my_sys_onchip_memory_s1_address),    //  output,   width = 7,                                                         my_sys_onchip_memory_s1.address
		.my_sys_onchip_memory_s1_write                                                         (mm_interconnect_0_my_sys_onchip_memory_s1_write),      //  output,   width = 1,                                                                                .write
		.my_sys_onchip_memory_s1_readdata                                                      (mm_interconnect_0_my_sys_onchip_memory_s1_readdata),   //   input,  width = 32,                                                                                .readdata
		.my_sys_onchip_memory_s1_writedata                                                     (mm_interconnect_0_my_sys_onchip_memory_s1_writedata),  //  output,  width = 32,                                                                                .writedata
		.my_sys_onchip_memory_s1_byteenable                                                    (mm_interconnect_0_my_sys_onchip_memory_s1_byteenable), //  output,   width = 4,                                                                                .byteenable
		.my_sys_onchip_memory_s1_chipselect                                                    (mm_interconnect_0_my_sys_onchip_memory_s1_chipselect), //  output,   width = 1,                                                                                .chipselect
		.my_sys_onchip_memory_s1_clken                                                         (mm_interconnect_0_my_sys_onchip_memory_s1_clken),      //  output,   width = 1,                                                                                .clken
		.mgc_axi4_master_0_reset_sink_reset_bridge_in_reset_reset                              (rst_controller_001_reset_out_reset),                   //   input,   width = 1,                              mgc_axi4_master_0_reset_sink_reset_bridge_in_reset.reset
		.mgc_axi4_master_0_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                   //   input,   width = 1, mgc_axi4_master_0_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset.reset
		.clock_in_out_clk_clk                                                                  (clock_in_out_clk_clk)                                  //   input,   width = 1,                                                                clock_in_out_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_in_out_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (clock_in_out_clk_clk),               //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (reset_in_out_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (clock_in_out_clk_clk),               //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
